class eth_mem_sequencer extends uvm_sequencer #(eth_sequence_item);

	`uvm_component_utils(eth_mem_sequencer)

	function new (string name="eth_mem_sequencer",uvm_component parent);
			super.new(name,parent);

	endfunction




endclass
